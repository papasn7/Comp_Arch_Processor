module rom_case(out, address);
	output reg [31:0] out;
	input  [31:0] address; // address- 16 deep memory  
	always @(address) begin
		case (address[31:2])
			16'h0000:  out = 32'b11010010100000000000000000100001; // MOVZ X1, 1
			16'h0001:  out = 32'b11010010100000000000000001000010; // MOVZ X2, 2
			16'h0002:  out = 32'b10001011000000100000000000100100; // ADD X4, X1, X2
			16'h0003:  out = 32'b11111000000000010000001111100100; // STUR X4, [XZR, 16]
			16'h0004:  out = 32'b11111000010000010000001111100101; // LDUR X5, [XZR, 16]
			16'h0005:  out = 32'b10010100000000000000000000001010; // BL 10
			16'h0006:  out = 32'b10110101000000000000000000100010; // CBNZ X2, 1
			16'h0007:  out = 32'b00010100000000000000000000000001; // B 1
			16'h0008:  out = 32'b00010111111111111111111111111001; // B -7
			16'h0009:  out = 32'b10110100000000000000000001100001; // CBZ X1, 3
			16'h000a:  out = 32'b11101011000000100000000000111111; // SUBS XZR, X1, X2
			16'h000b:  out = 32'b01010100000000000000000000100011; // B.LO 1
			16'h000c:  out = 32'b11111000000000001000001111100001; // STUR X1, [XZR, 8]
			16'h000d:  out = 32'b11111000010000001000001111100110; // LDUR X6, [XZR, 8]
			16'h000e:  out = 32'b11010010000000000000010011100111; // EORI X7, X7, 1
			16'h000f:  out = 32'b00010111111111111111111111111110; // B -2
			16'h0010:  out = 32'b10010001000000000000100000100001; // ADDI X1, X1, 2
			16'h0011:  out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
			16'h0012:  out = 32'b11010110000000000000001111000000; // BR X30
			default: out=32'b11010110000000000000000101100000; //BR X11
		endcase
	end
endmodule


/*
// Overclock (Nice!) Test
			// use X8 as the base address of RAM (default is 0x00000000)
			// For example if RAM is at 0x80000000 then change the following two instructions to:
			// MOVZ X8, 8 (put 8 in X8)
			// LSL X8, X8, 28 (shift it 28 times to get 0x80000000)
			16'h0000:  out = 32'b11010010100_0000000000000000_01000; // MOVZ X8, 0
			16'h0001:  out = 32'b1101001101100000_000000_0100001000; // LSL X8, X8, 0
			// use X11 as the base address of ROM (default is 0x00008000)
			16'h0002:  out = 32'b11010010100_0000000000001000_01011; // MOVZ X11, 8
			16'h0003:  out = 32'b1101001101100000_001100_0101101011; // LSL X11, X11, 12
			// X7 will hold the delay amount
			16'h0004:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 1
			// change the shift amount to change the delay
			// if using a testbench to debug then change the shift amount to 1
			16'h0005:  out = 32'b11010011011000000110000011100111; // LSL X7, X7, 24
			16'h0006:  out = 32'b11111000000000110000000100000111; // STUR X7, [X8, 48]
			16'h0007:  out = 32'b11010001000001100101011111100000; // SUBI X0, XZR, 405
			16'h0008:  out = 32'b11010001000100000000001111100101; // SUBI X5, XZR, 1024
			16'h0009:  out = 32'b10110010000001000110011111100010; // ORRI X2, XZR, 281
			16'h000a:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
			16'h000b:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
			16'h000c:  out = 32'b10001011000001010000000010100101; // ADD X5, X5, X5
			16'h000d:  out = 32'b10001011000000100000000010100010; // ADD X2, X5, X2
			16'h000e:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
			16'h000f:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
			16'h0010:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
			16'h0011:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
			16'h0012:  out = 32'b11001011000001010000001111100101; // SUB X5, XZR, X5
			16'h0013:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
			16'h0014:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
			16'h0015:  out = 32'b11111000000000011000000100000000; // STUR X0, [X8, 24]
			16'h0016:  out = 32'b11111000000000100000000100000010; // STUR X2, [X8, 32]
			16'h0017:  out = 32'b11111000000000101000000100000101; // STUR X5, [X8, 40]
			16'h0018:  out = 32'b10010001000000000000001111100000; // ADDI X0, XZR, 0
			16'h0019:  out = 32'b10010010000000000000001111100001; // ANDI X1, XZR, 0
			16'h001a:  out = 32'b11010010000000000000001111100010; // EORI X2, XZR, 0
			16'h001b:  out = 32'b10110010000000000000001111100011; // ORRI X3, XZR, 0
			16'h001c:  out = 32'b10101010000111110000001111100100; // ORR X4, X31, X31
			16'h001d:  out = 32'b10001010000111110000001111100101; // AND X5, X31, X31
			16'h001e:  out = 32'b10001010000111110000001111100110; // AND X6, X31, X31
			16'h001f:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
			16'h0020:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
			16'h0021:  out = 32'b10110101111111111111111111000111; // CBNZ X7, -2
			16'h0022:  out = 32'b11010010100111111111111111100000; // MOVZ X0, 65535
			16'h0023:  out = 32'b11010001000000000000011111100001; // SUBI X1, XZR, 1
			16'h0024:  out = 32'b11010010100111111111111111100010; // MOVZ X2, 65535
			16'h0025:  out = 32'b11010001000000000000011111100011; // SUBI X3, XZR, 1
			16'h0026:  out = 32'b11010010100111111111111111100100; // MOVZ X4, 65535
			16'h0027:  out = 32'b11010001000000000000011111100101; // SUBI X5, XZR, 1
			16'h0028:  out = 32'b11010001000000000000011111100110; // SUBI X6, XZR, 1
			16'h0029:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
			16'h002a:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
			16'h002b:  out = 32'b10110101111111111111111111000111; // CBNZ X7, -2
			16'h002c:  out = 32'b11111000010000011000000100000100; // LDUR X4, [X8, 24]
			16'h002d:  out = 32'b11111000010000100000000100000010; // LDUR X2, [X8, 32]
			16'h002e:  out = 32'b11111000010000101000000100000101; // LDUR X5, [X8, 40]
			16'h002f:  out = 32'b10010001000000000000000001000011; // ADDI X3, X2, 0
			16'h0030:  out = 32'b10110010000000010000000001100011; // ORRI X3, X3, 64
			16'h0031:  out = 32'b11010010100000000000000100000111; // MOVZ X7, 8
			16'h0032:  out = 32'b11001011000001110000000001100011; // SUB X3, X3, X7
			16'h0033:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 1
			16'h0034:  out = 32'b11001010000001110000000001100001; // EOR X1, X3, X7
			16'h0035:  out = 32'b11001011000001010000000000100001; // SUB X1, X1, X5
			16'h0036:  out = 32'b10110010000000000000000010000000; // ORRI X0, X4, 0
			16'h0037:  out = 32'b11010010100000000000000000000101; // MOVZ X5, 0
			16'h0038:  out = 32'b11010010100000000000000000000110; // MOVZ X6, 0
			16'h0039:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
			16'h003a:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
			16'h003b:  out = 32'b10110101111111111111111111000111; // CBNZ X7, -2
			16'h003c:  out = 32'b11010110000000000000000101100000; // BR X11
			default: out=32'b11010110000000000000000101100000; //BR X11
*/

/*			ECE
			16'h0000:  out = 32'b11010010100111110011101111100000; // MOVZ X0, 63967
			16'h0001:  out = 32'b11010010100000000000000000101010; // MOVZ X10, 1
			16'h0002:  out = 32'b11010011011000000010100101001010; // LSL X10, X10, 10
			16'h0003:  out = 32'b11111000000000000000000101000000; // STUR X0, [X10, 0]																		 // 
			16'h0004:  out = 32'b11010010100100000100001000000001; // MOVZ X1, 33296
			16'h0005:  out = 32'b11010010100000000000000000101011; // MOVZ X11, 1
			16'h0006:  out = 32'b11010011011000000010110101101011; // LSL X11, X11, 11
			16'h0007:  out = 32'b11111000000000000000000101100001; // STUR X1, [X11, 0]
			16'h0008:  out = 32'b11010010100100000100001000000010; // MOVZ X2, 33296
			16'h0009:  out = 32'b11010010100000000000000000101100; // MOVZ X12, 1
			16'h000a:  out = 32'b11010011011000000011000110001100; // LSL X12, X12, 12
			16'h000b:  out = 32'b11111000000000000000000110000010; // STUR X2, [X12, 0]
			16'h000c:  out = 32'b11010010100100000100001000000011; // MOVZ X3, 33296
			16'h000d:  out = 32'b11010010100000000000000000101101; // MOVZ X13, 1
			16'h000e:  out = 32'b11010011011000000011010110101101; // LSL X13, X13, 13
			16'h000f:  out = 32'b11111000000000000000000110100011; // STUR X3, [X13, 0]
			16'h0010:  out = 32'b11010010100111100100001111000100; // MOVZ X4, 61982
			16'h0011:  out = 32'b11010010100000000000000000101110; // MOVZ X14, 1
			16'h0012:  out = 32'b11010011011000000011100111001110; // LSL X14, X14, 14
			16'h0013:  out = 32'b11111000000000000000000111000100; // STUR X4, [X14, 0]
			16'h0014:  out = 32'b11010010100100000100001000000101; // MOVZ X5, 33296
			16'h0015:  out = 32'b11010010100000000000000000101111; // MOVZ X15, 1
			16'h0016:  out = 32'b11010011011000000011110111101111; // LSL X15, X15, 15
			16'h0017:  out = 32'b11111000000000000000000111100101; // STUR X5, [X15, 0]
			16'h0018:  out = 32'b11010010100100000100001000000110; // MOVZ X6, 33296
			16'h0019:  out = 32'b11010010100000000000000000110000; // MOVZ X16, 1
			16'h001a:  out = 32'b11010011011000000100001000010000; // LSL X16, X16, 16
			16'h001b:  out = 32'b11111000000000000000001000000110; // STUR X6, [X16, 0]
			16'h001c:  out = 32'b11010010100111110011101111100111; // MOVZ X7, 63967
			16'h001d:  out = 32'b11010010100000000000000000110001; // MOVZ X17, 1
			16'h001e:  out = 32'b11010011011000000100011000110001; // LSL X17, X17, 17
			16'h001f:  out = 32'b11111000000000000000001000100111; // STUR X7, [X17, 0]
*/

/*
			16'h0000:  out = 32'b11010010100111110010000111000000; // MOVZ X0, 63758
			16'h0001:  out = 32'b11010010100000000000000000101010; // MOVZ X10, 1
			16'h0002:  out = 32'b11010011011000000010100101001010; // LSL X10, X10, 10
			16'h0003:  out = 32'b11010010100001000010001000100001; // MOVZ X1, 8465
			16'h0004:  out = 32'b11010010100000000000000000101011; // MOVZ X11, 1
			16'h0005:  out = 32'b11010011011000000010110101101011; // LSL X11, X11, 11
			16'h0006:  out = 32'b11010010100001000101001000100010; // MOVZ X2, 8849
			16'h0007:  out = 32'b11010010100000000000000000101100; // MOVZ X12, 1
			16'h0008:  out = 32'b11010011011000000011000110001100; // LSL X12, X12, 12
			16'h0009:  out = 32'b11010010100001001000101000100011; // MOVZ X3, 9297
			16'h000a:  out = 32'b11010010100000000000000000101101; // MOVZ X13, 1
			16'h000b:  out = 32'b11010011011000000011010110101101; // LSL X13, X13, 13
			16'h000c:  out = 32'b11010010100001010000011000100100; // MOVZ X4, 10289
			16'h000d:  out = 32'b11010010100000000000000000101110; // MOVZ X14, 1
			16'h000e:  out = 32'b11010011011000000011100111001110; // LSL X14, X14, 14
			16'h000f:  out = 32'b11010010100001010010011000100101; // MOVZ X5, 10545
			16'h0010:  out = 32'b11010010100000000000000000101111; // MOVZ X15, 1
			16'h0011:  out = 32'b11010011011000000011110111101111; // LSL X15, X15, 15
			16'h0012:  out = 32'b11010010100001001101101000100110; // MOVZ X6, 9937
			16'h0013:  out = 32'b11010010100000000000000000110000; // MOVZ X16, 1
			16'h0014:  out = 32'b11010011011000000100001000010000; // LSL X16, X16, 16
			16'h0015:  out = 32'b11010010100111110000001000100111; // MOVZ X7, 63505
			16'h0016:  out = 32'b11010010100000000000000000110001; // MOVZ X17, 1
			16'h0017:  out = 32'b11010011011000000100011000110001; // LSL X17, X17, 17
*/